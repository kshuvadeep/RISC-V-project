// Memory control macros
`define CTRL_MEM_WIDTH 3 
`define CTRL_LB  3'b000  // Load Byte
`define CTRL_LH  3'b001  // Load Halfword
`define CTRL_LW  3'b010  // Load Word
`define CTRL_LBU 3'b011  // Load Byte Unsigned
`define CTRL_LHU 3'b100  // Load Halfword Unsigned

`define CTRL_SB  3'b000  // Store Byte
`define CTRL_SH  3'b001  // Store Halfword
`define CTRL_SW  3'b010  // Store Word
