//*******************
//this file  contains the crucial 
//system parameter like address width ,data width , 
//and other such parameters 

`define DATA_WIDTH 32 
`define ADDR_WIDTH 32 
