
// defines for adder
`define CTRL_ADD_WIDTH 2 
`define CTRL_ADD 2'b01
`define CTRL_SUB 2'b10
`define CTRL_ADDI 2'b11

//defines for shifter 


//defines for logic 
`define CTRL_LOGIC_WIDTH 3
`define CTRL_XOR 3'b000
`define CTRL_OR 3'b001
`define CTRL_AND 3'b010
`define CTRL_ANDI 3'b101
`define CTRL_XORI 3'b111
`define CTRL_ORI 3'b110
`define MSB_CTRL 2

