//*******************
//this file  contains the crucial 
//system parameter like address width ,data width , 
//and other such parameters 


`define DATA_WIDTH 32 
`define DATA_WIDTH 32 
`define INST_WIDTH 32 
`define REG_ADDR_WIDTH 5  
`define ADDR_WIDTH 32
`define OPCODE_WIDTH 7 
`define IMMEDIATE_WIDTH 21
`define MEM_DATA_WIDTH 8
`define IO_SELECT 4 
`define MEM_DEPTH 64 
//CSN SELECT

`define MEM_SELECT 4'b0000
`define UART_SELECT 4'b1000 
