
// defines for adder 
`define CTRL_ADD 2'b01
`define CTRL_SUB 2'b10
`define CTRL_ADDI 2'b11

//defines for shifter 

