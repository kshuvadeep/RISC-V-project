
`define zero 5'b00000   // Hardwired zero
`define ra   5'b00001   // Return address
`define sp   5'b00010   // Stack pointer
`define gp   5'b00011   // Global pointer
`define tp   5'b00100   // Thread pointer
`define t0   5'b00101   // Temporary
`define t1   5'b00110   // Temporary
`define t2   5'b00111   // Temporary
`define s0   5'b01000   // Saved register/frame pointer
`define fp   5'b01000   // Frame pointer (alias for s0)
`define s1   5'b01001   // Saved register
`define a0   5'b01010   // Function argument/return value
`define a1   5'b01011   // Function argument/return value
`define a2   5'b01100   // Function argument
`define a3   5'b01101   // Function argument
`define a4   5'b01110   // Function argument
`define a5   5'b01111   // Function argument
`define a6   5'b10000   // Function argument
`define a7   5'b10001   // Function argument
`define s2   5'b10010   // Saved register
`define s3   5'b10011   // Saved register
`define s4   5'b10100   // Saved register
`define s5   5'b10101   // Saved register
`define s6   5'b10110   // Saved register
`define s7   5'b10111   // Saved register
`define s8   5'b11000   // Saved register
`define s9   5'b11001   // Saved register
`define s10  5'b11010   // Saved register
`define s11  5'b11011   // Saved register
`define t3   5'b11100   // Temporary
`define t4   5'b11101   // Temporary
`define t5   5'b11110   // Temporary
`define t6   5'b11111   // Temporary
