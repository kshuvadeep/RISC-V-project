// This module consists of UArt tx , uart rx ,and Fifo .
// This module works as an IO module connected to main
// cpu core via a system bus .
//We will use Memory mapped IO to send data to it
//Uart works as an interface to send data to any other devices
//It can be a raspberry pi or a laptop
// Author: Shuvadeep Kumar

//Date :22nd october

`include "system_param.vh"
`include "Macros.vh"

module Uart_module(
         input clk ,
         input reset,
         //system bus
         input[`ADDR_WIDTH-1:0] addr ,
         inout[`DATA_WIDTH-1:0] wrt_data ,
         output[`DATA_WIDTH-1:0] rd_data ,
         input programming,
         input we ,
         input req_valid,
         output data_valid ,   // will work as ready for read operation
         //
         output txd ,
         input rxd
       );

       wire packet_v;
      wire [`DATA_WIDTH-1:0] data_packet;
      wire [`DATA_WIDTH-1:0] rd_data_rx;


      reg wrt_clk_tx;
      wire rd_clk_tx;
      reg wrt_clk_rx, rd_clk_rx;
      wire [`DATA_WIDTH-1:0] tx_data;
     //subscript tx and rx stands for the corresponding modules
      wire wrt_en_tx ,rd_en_tx;
      wire wrt_en_rx, rd_en_rx ;
      wire tx_enable ,rx_enable  ;
      wire tx_full , tx_empty ;
      wire csn_uart ; // whether the Uart module is selected or not
      wire Uart_out_valid ;
      wire[7:0] Uart_data_out;
      wire data_valid_arbiter;

       // chip select login
       assign csn_uart =  (addr[`ADDR_WIDTH-1: `ADDR_WIDTH-`IO_SELECT] ==`UART_SELECT ) ? 1'b1 :1'b0;

      //rd and wrt enbale logic
      assign wrt_en_tx = req_valid & csn_uart & we ;
      assign rd_en_tx = !tx_empty & tx_enable ;


   //   assign rd_en_rx <= req_valid & (addr[`ADDR_WIDTH: `ADDR_WIDTH-`IO_SELECT] ==4'b0001 ) & !we ;
   //   assign wrt_en_rx <= !rx_empty & rx_enable  ;

     // `CLK_GATE(clk,wrt_en_tx,wrt_clk_tx)
    always@(*) begin
     wrt_clk_tx =  wrt_en_tx;
   end
     // `CLK_GATE(clk,rd_en_tx,rd_clk_tx)

   //   CLK_GATE(clk,wrt_en_rx,wrt_clk_rx)
   //   CLK_GATE(clk,rd_en_rx,rd_clk_rx)


      //Fifo for TX

       Fifo #(
        .DEPTH(16),      // Set depth of FIFO to 16
        .WIDTH(32)       // Set width of data to 32 bits
    ) fifo_tx (
        .reset(reset),
        .wrt_clk(wrt_clk_tx),
        .rd_clk(rd_clk_tx),
        .wrt_data(wrt_data),
        .rd_data(tx_data),
        .full(tx_full),
        .empty(tx_empty)
    );



     // Transmission module

   Uart_tx uart_tx_inst (
        .clk(clk),
        .reset(reset),
        .data(tx_data),
        .tx_fifo_empty(tx_empty),
        .rd_clk_tx(rd_clk_tx),
        .txd(txd)
    );

     //receiving module ,currently just testing the functionality

  Uart_rx  #(.CLK_FREQ(50) , .BAUD_RATE(9600))
       Uart_rx_inst     (
     .i_clk(clk),
     .i_Rx_Serial(rxd) ,
     .o_Rx_DV(Uart_out_valid),
     .o_Rx_Byte(Uart_data_out)
     );


  packet_builder #( .NUM_BYTE(4))
      uart_packet_builder
        (
                .clk(clk),
                 .rst(reset),
                .data_byte(Uart_data_out),
                .data_byte_valid(Uart_out_valid),
                .packet_data(data_packet),
                .packet_valid(packet_v)
        );

   Arbiter_uart_rx
     u_Arbiter_uart_rx (
      .clk(clk),
      .rst(reset),
      //address
      .addr(addr),
      //data
      .packet_v(packet_v),
      .packet_data(data_packet),
      .wrt_data(wrt_data),
      .rd_data(rd_data_rx),
      //control signals
      .programming(programming),
      .csn_uart(csn_uart),
       // output ready ,// optional ,to tell the sender it's status .
     .req_valid(req_valid),
     .data_valid(data_valid),
     .arbiter_data_valid(data_valid_arbiter),
     .we(we)
 );



     assign data_valid = programming ? 1'bz : csn_uart ? (!tx_full| data_valid_arbiter  ):1'bz; // needs to  modify this for the Receiver module

   // since the RX module is not designed yet
    assign rd_data = csn_uart ? rd_data_rx : {`DATA_WIDTH{1'bz}};


endmodule
